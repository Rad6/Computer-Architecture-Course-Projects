library verilog;
use verilog.vl_types.all;
entity HazardDetecting_TB is
end HazardDetecting_TB;
