library verilog;
use verilog.vl_types.all;
entity Controller is
    generic(
        \IF\            : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        ID              : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        JMP1            : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi1, Hi0);
        JZ1             : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi1, Hi1);
        PUSH1           : vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi0, Hi0);
        PUSH2           : vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi0, Hi1);
        O1              : vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi1, Hi0);
        O2              : vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi1, Hi1);
        POP1            : vl_logic_vector(3 downto 0) := (Hi1, Hi0, Hi0, Hi0);
        NOT1            : vl_logic_vector(3 downto 0) := (Hi1, Hi0, Hi0, Hi1);
        PUSHG           : vl_logic_vector(3 downto 0) := (Hi1, Hi0, Hi1, Hi0);
        LOGIC1          : vl_logic_vector(3 downto 0) := (Hi1, Hi0, Hi1, Hi1);
        LOGIC2          : vl_logic_vector(3 downto 0) := (Hi1, Hi1, Hi0, Hi0);
        LOGIC3          : vl_logic_vector(3 downto 0) := (Hi1, Hi1, Hi0, Hi1);
        \_push\         : vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        \_pop\          : vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi1);
        \_jmp\          : vl_logic_vector(2 downto 0) := (Hi1, Hi1, Hi0);
        \_jz\           : vl_logic_vector(2 downto 0) := (Hi1, Hi1, Hi1);
        \_add\          : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        \_sub\          : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi1);
        \_and\          : vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi0);
        \_not\          : vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi1);
        alu_sub         : vl_logic_vector(1 downto 0) := (Hi0, Hi1);
        alu_add         : vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        alu_and         : vl_logic_vector(1 downto 0) := (Hi1, Hi0);
        alu_not         : vl_logic_vector(1 downto 0) := (Hi1, Hi1)
    );
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        inst            : in     vl_logic_vector(2 downto 0);
        PcWrite         : out    vl_logic;
        PcWriteC        : out    vl_logic;
        PcSrc           : out    vl_logic;
        PorI            : out    vl_logic;
        MemRead         : out    vl_logic;
        IRWrite         : out    vl_logic;
        MemWrite        : out    vl_logic;
        MtoS            : out    vl_logic;
        LdA             : out    vl_logic;
        LdB             : out    vl_logic;
        SrcA            : out    vl_logic;
        SrcB            : out    vl_logic;
        Push            : out    vl_logic;
        Pop             : out    vl_logic;
        toS             : out    vl_logic;
        AluOp           : out    vl_logic_vector(1 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of \IF\ : constant is 2;
    attribute mti_svvh_generic_type of ID : constant is 2;
    attribute mti_svvh_generic_type of JMP1 : constant is 2;
    attribute mti_svvh_generic_type of JZ1 : constant is 2;
    attribute mti_svvh_generic_type of PUSH1 : constant is 2;
    attribute mti_svvh_generic_type of PUSH2 : constant is 2;
    attribute mti_svvh_generic_type of O1 : constant is 2;
    attribute mti_svvh_generic_type of O2 : constant is 2;
    attribute mti_svvh_generic_type of POP1 : constant is 2;
    attribute mti_svvh_generic_type of NOT1 : constant is 2;
    attribute mti_svvh_generic_type of PUSHG : constant is 2;
    attribute mti_svvh_generic_type of LOGIC1 : constant is 2;
    attribute mti_svvh_generic_type of LOGIC2 : constant is 2;
    attribute mti_svvh_generic_type of LOGIC3 : constant is 2;
    attribute mti_svvh_generic_type of \_push\ : constant is 2;
    attribute mti_svvh_generic_type of \_pop\ : constant is 2;
    attribute mti_svvh_generic_type of \_jmp\ : constant is 2;
    attribute mti_svvh_generic_type of \_jz\ : constant is 2;
    attribute mti_svvh_generic_type of \_add\ : constant is 2;
    attribute mti_svvh_generic_type of \_sub\ : constant is 2;
    attribute mti_svvh_generic_type of \_and\ : constant is 2;
    attribute mti_svvh_generic_type of \_not\ : constant is 2;
    attribute mti_svvh_generic_type of alu_sub : constant is 2;
    attribute mti_svvh_generic_type of alu_add : constant is 2;
    attribute mti_svvh_generic_type of alu_and : constant is 2;
    attribute mti_svvh_generic_type of alu_not : constant is 2;
end Controller;
