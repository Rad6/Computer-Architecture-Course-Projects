library verilog;
use verilog.vl_types.all;
entity stack_TB is
end stack_TB;
