library verilog;
use verilog.vl_types.all;
entity IM_TB is
end IM_TB;
