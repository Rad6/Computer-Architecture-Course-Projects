library verilog;
use verilog.vl_types.all;
entity TB_IfZero is
end TB_IfZero;
