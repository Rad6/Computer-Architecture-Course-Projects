library verilog;
use verilog.vl_types.all;
entity TB_RF is
end TB_RF;
