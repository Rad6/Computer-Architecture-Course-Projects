library verilog;
use verilog.vl_types.all;
entity TB_PIPELINE is
end TB_PIPELINE;
