library verilog;
use verilog.vl_types.all;
entity TB_ForwardingUnit is
end TB_ForwardingUnit;
