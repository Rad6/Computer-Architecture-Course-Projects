library verilog;
use verilog.vl_types.all;
entity FILEREADER_TB is
end FILEREADER_TB;
