library verilog;
use verilog.vl_types.all;
entity TB_MIPS is
end TB_MIPS;
