module ROM(input [7:0] address, output reg signed [15:0] data);
  always @(address)
  case (address)
    0  : data = 16'b0001101000100101;
    1  : data = 16'b0010010001100001;
    2  : data = 16'b0010010001000001;
    3  : data = 16'b0000010001101101;
    4  : data = 16'b0000110000011101;
    5  : data = 16'b0000010001001001;
    6  : data = 16'b0001111000100001;
    7  : data = 16'b0000010001010101;
    8  : data = 16'b0010110001101001;
    9  : data = 16'b0001000001100001;
    10 : data = 16'b0000111111111101;
    11 : data = 16'b0011110001010101;
    12 : data = 16'b0100001001000001;
    13 : data = 16'b0001001001001101;
    14 : data = 16'b0010000000110001;
    15 : data = 16'b0100000000001101;
    16 : data = 16'b0001100001011101;
    17 : data = 16'b0011110000110001;
    18 : data = 16'b0010111000110101;
    19 : data = 16'b0010000001000101;
    20 : data = 16'b0001101010010001;
    21 : data = 16'b0011110010001001;
    22 : data = 16'b0010110000010101;
    23 : data = 16'b0001011000110001;
    24 : data = 16'b0010011001100001;
    25 : data = 16'b0001001111111101;
    26 : data = 16'b0010001001101001;
    27 : data = 16'b0011100000110101;
    28 : data = 16'b0010100001101101;
    29 : data = 16'b0001010000100101;
    30 : data = 16'b0010011000100101;
    31 : data = 16'b0001010010001101;
    32 : data = 16'b0100000001010101;
    33 : data = 16'b0000010000111001;
    34 : data = 16'b0001011000100001;
    35 : data = 16'b0010110001100101;
    36 : data = 16'b0001001001001101;
    37 : data = 16'b0010000111111001;
    38 : data = 16'b0010101000100101;
    39 : data = 16'b0011010010100001;
    40 : data = 16'b0001001001000001;
    41 : data = 16'b0001111000000001;
    42 : data = 16'b0001100000100101;
    43 : data = 16'b0001111000110101;
    44 : data = 16'b0010011001011001;
    45 : data = 16'b0001011000111101;
    46 : data = 16'b0010110001000101;
    47 : data = 16'b0010011001000001;
    48 : data = 16'b0001100000100001;
    49 : data = 16'b0010010001100101;
    50 : data = 16'b0011000000110101;
    51 : data = 16'b0011000000110001;
    52 : data = 16'b0010101001001001;
    53 : data = 16'b0001111000111101;
    54 : data = 16'b0001011000110001;
    55 : data = 16'b0010010001000101;
    56 : data = 16'b0001100010000101;
    57 : data = 16'b0001101001010001;
    58 : data = 16'b0010111000101101;
    59 : data = 16'b0011100000100101;
    60 : data = 16'b0010101000111001;
    61 : data = 16'b0100000000001101;
    62 : data = 16'b0000100001111101;
    63 : data = 16'b0010000001001001;
    64 : data = 16'b0010001000011101;
    65 : data = 16'b0011101001000101;
    66 : data = 16'b0010100000010001;
    67 : data = 16'b0001101001010101;
    68 : data = 16'b0010100000111101;
    69 : data = 16'b0010101001000001;
    70 : data = 16'b0010001001001101;
    71 : data = 16'b0000000001011101;
    72 : data = 16'b0011000000101001;
    73 : data = 16'b1110100000010001;
    74 : data = 16'b0010001000111101;
    75 : data = 16'b0000100000100101;
    76 : data = 16'b0001101001001101;
    77 : data = 16'b0011011000000101;
    78 : data = 16'b0001100001011101;
    79 : data = 16'b0011111001001001;
    80 : data = 16'b0010110000011101;
    81 : data = 16'b0001110000110101;
    82 : data = 16'b0001001001011101;
    83 : data = 16'b0001100010001101;
    84 : data = 16'b0010011000110101;
    85 : data = 16'b1111101001101101;
    86 : data = 16'b0010101000100101;
    87 : data = 16'b0010010001001001;
    88 : data = 16'b0010111000111001;
    89 : data = 16'b0100000001001101;
    90 : data = 16'b0001101000110001;
    91 : data = 16'b0001000000010101;
    92 : data = 16'b0011001000111001;
    93 : data = 16'b0010111001010001;
    94 : data = 16'b0001111000110001;
    95 : data = 16'b0001011000111101;
    96 : data = 16'b0010010001001101;
    97 : data = 16'b0000111001010001;
    98 : data = 16'b0010001000101001;
    99 : data = 16'b0001011000111001;
    100: data = 16'b1110111110101011;
    101: data = 16'b1110011110100111;
    102: data = 16'b1100101111111011;
    103: data = 16'b1111100110100111;
    104: data = 16'b1101011110111011;
    105: data = 16'b1101010110100111;
    106: data = 16'b1100101111011111;
    107: data = 16'b1101111111000011;
    108: data = 16'b1101111111000111;
    109: data = 16'b1101101111100011;
    110: data = 16'b1101001111010111;
    111: data = 16'b1100011111011011;
    112: data = 16'b0001000101111111;
    113: data = 16'b1111100111001011;
    114: data = 16'b1101101111100011;
    115: data = 16'b1101111111001111;
    116: data = 16'b1110011111011111;
    117: data = 16'b1110000000000111;
    118: data = 16'b1101011111101011;
    119: data = 16'b1110111110011111;
    120: data = 16'b1100111110100111;
    121: data = 16'b0000000110111111;
    122: data = 16'b1100010110101111;
    123: data = 16'b1101101110111111;
    124: data = 16'b1110111111101011;
    125: data = 16'b1110001110110011;
    126: data = 16'b1100100110111011;
    127: data = 16'b1110111110111011;
    128: data = 16'b1110001111010111;
    129: data = 16'b1101001111100011;
    130: data = 16'b1110011110111111;
    131: data = 16'b1110110110110111;
    132: data = 16'b0000001111011111;
    133: data = 16'b1101111111011011;
    134: data = 16'b1101110111010011;
    135: data = 16'b1101100000101011;
    136: data = 16'b1100001111000011;
    137: data = 16'b1110100111001111;
    138: data = 16'b1100000110111111;
    139: data = 16'b1101110111010111;
    140: data = 16'b1101110110110011;
    141: data = 16'b1110111111100011;
    142: data = 16'b1011010111111111;
    143: data = 16'b1110111111000111;
    144: data = 16'b1101100110111111;
    145: data = 16'b1100110110101111;
    146: data = 16'b1110000110110011;
    147: data = 16'b1110010110001011;
    148: data = 16'b1101101111000011;
    149: data = 16'b1100100110100111;
    150: data = 16'b1111010111101011;
    151: data = 16'b1110010111000111;
    152: data = 16'b1101010111000011;
    153: data = 16'b1111010111101111;
    154: data = 16'b1110011110001011;
    155: data = 16'b1100110111001111;
    156: data = 16'b1110101110100011;
    157: data = 16'b1100010110101111;
    158: data = 16'b1101000111001011;
    159: data = 16'b1110001111011111;
    160: data = 16'b1110011110100111;
    161: data = 16'b1110001111010011;
    162: data = 16'b1100001111110011;
    163: data = 16'b1110111110100111;
    164: data = 16'b1111010110100011;
    165: data = 16'b1111001111000011;
    166: data = 16'b1101011111010111;
    167: data = 16'b1101101111000011;
    168: data = 16'b1101000110100111;
    169: data = 16'b1110010111000111;
    170: data = 16'b1110010111001011;
    171: data = 16'b1101010110110011;
    172: data = 16'b1110111110011111;
    173: data = 16'b1110111111001111;
    174: data = 16'b1110101111000011;
    175: data = 16'b1101010110110111;
    176: data = 16'b1100101110101111;
    177: data = 16'b1110101110110011;
    178: data = 16'b1111100110100111;
    179: data = 16'b1100110110100011;
    180: data = 16'b1011110111101011;
    181: data = 16'b1111011110111011;
    182: data = 16'b1110000110001011;
    183: data = 16'b1111001110110011;
    184: data = 16'b1111000111100011;
    185: data = 16'b1100110110110011;
    186: data = 16'b1101101111111011;
    187: data = 16'b1101001110101011;
    188: data = 16'b1110001110101011;
    189: data = 16'b1111001110100011;
    190: data = 16'b1110000111100111;
    191: data = 16'b1011111110101111;
    192: data = 16'b1111010111001111;
    193: data = 16'b1110000110001111;
    194: data = 16'b1101100110101111;
    195: data = 16'b1011111111010111;
    196: data = 16'b1110011110011011;
    197: data = 16'b1110010111000011;
    198: data = 16'b1110011111010011;
    199: data = 16'b1100111111111011;
  endcase
endmodule







// list = ['0001101000100101',
//   '0010010001000001',
//   '0010010001100001',
//   '0000010001101101',
//   '0000110000011101',
//   '0000010001001001',
//   '0001111000100001',
//   '0000010001010101',
//   '0010110001101001',
//   '0001000001100001',
//   '0000111111111101',
//   '0011110001010101',
//   '0100001001000001',
//   '0001001001001101',
//   '0010000000110001',
//   '0100000000001101',
//   '0001100001011101',
//   '0011110000110001',
//   '0010111000110101',
//   '0010000001000101',
//   '0001101010010001',
//   '0011110010001001',
//   '0010110000010101',
//   '0001011000110001',
//   '0010011001100001',
//   '0001001111111101',
//   '0010001001101001',
//   '0011100000110101',
//   '0010100001101101',
//   '0001010000100101',
//   '0010011000100101',
//   '0001010010001101',
//   '0100000001010101',
//   '0000010000111001',
//   '0001011000100001',
//   '0010110001100101',
//   '0001001001001101',
//   '0010000111111001',
//   '0010101000100101',
//   '0011010010100001',
//   '0001001001000001',
//   '0001111000000001',
//   '0001100000100101',
//   '0001111000110101',
//   '0010011001011001',
//   '0001011000111101',
//   '0010110001000101',
//   '0010011001000001',
//   '0001100000100001',
//   '0010010001100101',
//   '0011000000110101',
//   '0011000000110001',
//   '0010101001001001',
//   '0001111000111101',
//   '0001011000110001',
//   '0010010001000101',
//   '0001100010000101',
//   '0001101001010001',
//   '0010111000101101',
//   '0011100000100101',
//   '0010101000111001',
//   '0100000000001101',
//   '0000100001111101',
//   '0010000001001001',
//   '0010001000011101',
//   '0011101001000101',
//   '0010100000010001',
//   '0001101001010101',
//   '0010100000111101',
//   '0010101001000001',
//   '0010001001001101',
//   '0000000001011101',
//   '0011000000101001',
//   '1110100000010001',
//   '0010001000111101',
//   '0000100000100101',
//   '0001101001001101',
//   '0011011000000101',
//   '0001100001011101',
//   '0011111001001001',
//   '0010110000011101',
//   '0001110000110101',
//   '0001001001011101',
//   '0001100010001101',
//   '0010011000110101',
//   '1111101001101101',
//   '0010101000100101',
//   '0010010001001001',
//   '0010111000111001',
//   '0100000001001101',
//   '0001101000110001',
//   '0001000000010101',
//   '0011001000111001',
//   '0010111001010001',
//   '0001111000110001',
//   '0001011000111101',
//   '0010010001001101',
//   '0000111001010001',
//   '0010001000101001',
//   '0001011000111001',
//   '1110111110101011',
//   '1110011110100111',
//   '1100101111111011',
//   '1111100110100111',
//   '1101011110111011',
//   '1101010110100111',
//   '1100101111011111',
//   '1101111111000011',
//   '1101111111000111',
//   '1101101111100011',
//   '1101001111010111',
//   '1100011111011011',
//   '0001000101111111',
//   '1111100111001011',
//   '1101101111100011',
//   '1101111111001111',
//   '1110011111011111',
//   '1110000000000111',
//   '1101011111101011',
//   '1110111110011111',
//   '1100111110100111',
//   '0000000110111111',
//   '1100010110101111',
//   '1101101110111111',
//   '1110111111101011',
//   '1110001110110011',
//   '1100100110111011',
//   '1110111110111011',
//   '1110001111010111',
//   '1101001111100011',
//   '1110011110111111',
//   '1110110110110111',
//   '0000001111011111',
//   '1101111111011011',
//   '1101110111010011',
//   '1101100000101011',
//   '1100001111000011',
//   '1110100111001111',
//   '1100000110111111',
//   '1101110111010111',
//   '1101110110110011',
//   '1110111111100011',
//   '1011010111111111',
//   '1110111111000111',
//   '1101100110111111',
//   '1100110110101111',
//   '1110000110110011',
//   '1110010110001011',
//   '1101101111000011',
//   '1100100110100111',
//   '1111010111101011',
//   '1110010111000111',
//   '1101010111000011',
//   '1111010111101111',
//   '1110011110001011',
//   '1100110111001111',
//   '1110101110100011',
//   '1100010110101111',
//   '1101000111001011',
//   '1110001111011111',
//   '1110011110100111',
//   '1110001111010011',
//   '1100001111110011',
//   '1110111110100111',
//   '1111010110100011',
//   '1111001111000011',
//   '1101011111010111',
//   '1101101111000011',
//   '1101000110100111',
//   '1110010111000111',
//   '1110010111001011',
//   '1101010110110011',
//   '1110111110011111',
//   '1110111111001111',
//   '1110101111000011',
//   '1101010110110111',
//   '1100101110101111',
//   '1110101110110011',
//   '1111100110100111',
//   '1100110110100011',
//   '1011110111101011',
//   '1111011110111011',
//   '1110000110001011',
//   '1111001110110011',
//   '1111000111100011',
//   '1100110110110011',
//   '1101101111111011',
//   '1101001110101011',
//   '1110001110101011',
//   '1111001110100011',
//   '1110000111100111',
//   '1011111110101111',
//   '1111010111001111',
//   '1110000110001111',
//   '1101100110101111',
//   '1011111111010111',
//   '1110011110011011',
//   '1110010111000011',
//   '1110011111010011',
//   '1100111111111011']


// for i in range(len(list)):
//   print(int(list[i],2))