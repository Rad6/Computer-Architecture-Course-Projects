library verilog;
use verilog.vl_types.all;
entity TB_MEM is
end TB_MEM;
