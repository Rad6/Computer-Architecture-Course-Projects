library verilog;
use verilog.vl_types.all;
entity PC_TB is
end PC_TB;
