library verilog;
use verilog.vl_types.all;
entity RegFile_TB is
end RegFile_TB;
