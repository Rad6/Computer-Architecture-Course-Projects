library verilog;
use verilog.vl_types.all;
entity MEM_TB is
end MEM_TB;
