library verilog;
use verilog.vl_types.all;
entity cache_tb is
end cache_tb;
